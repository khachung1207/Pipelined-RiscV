module And_module(
	 input logic [31:0] And_A, And_B,
	 output logic [31:0] And_kq
);

assign And_kq = And_A & And_B; 
endmodule 